library verilog;
use verilog.vl_types.all;
entity convert2Disp7_vlg_vec_tst is
end convert2Disp7_vlg_vec_tst;
