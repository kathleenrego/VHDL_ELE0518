library verilog;
use verilog.vl_types.all;
entity convert3Disp_vlg_vec_tst is
end convert3Disp_vlg_vec_tst;
