library verilog;
use verilog.vl_types.all;
entity Lab7_vlg_vec_tst is
end Lab7_vlg_vec_tst;
